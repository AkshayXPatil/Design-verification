interface ram_intf (input logic clk,rst);

logic [3:0] addr, idata, odata;
logic wr,en;

endinterface